dfdjk
